module 400g_axis_adapter #(
    parameter ETH = 400
)(

);

endmodule