module 400g_axis_adapter_sim;

endmodule;